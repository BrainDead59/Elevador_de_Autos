library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.std_logic_arith.ALL;
use IEEE.std_logic_unsigned.ALL;

entity DivisorServomotor is
	port(clk: in std_logic;
		  div_clk: out std_logic);
end DivisorServomotor;

architecture Behavioral of DivisorServomotor is
begin
	process(clk)
		constant N: integer :=3;
		variable cuenta: std_logic_vector(27 downto 0) :=X"0000000";
	begin
		if rising_edge(clk) then
			cuenta:=cuenta+1;
		end if;
		div_clk <= cuenta(N);
	end process;
end Behavioral;
